`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/30/2024 12:12:06 PM
// Design Name: 
// Module Name: tb_Encryption
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module tb_Decryption;

  // Parameters
  parameter N = 3;
  parameter d = 4;

  // Signals
    reg clk;
    reg reset;
    reg [N-1:0] x_C1;
    reg [N-1:0] y_C1;
    reg [N-1:0] z_C1;
    reg [N-1:0] x_C2;
    reg [N-1:0] y_C2;
    reg [N-1:0] z_C2;
    wire [N-1:0] x_Plaintext;
    wire [N-1:0] y_Plaintext;
    wire [N-1:0] z_Plaintext;
    wire Decryption_ready;
  // Instantiate the module under test
  Decryption #(
        .N(N),
        .ds(d)
       
  ) dut (
    .clk(clk),
    .reset(reset),
    .x_C1(x_C1),
    .y_C1(y_C1),
    .z_C1(z_C1),
    .x_C2(x_C2),
    .y_C2(y_C2),
    .z_C2(z_C2),
    .x_Plaintext(x_Plaintext),
    .y_Plaintext(y_Plaintext),
    .z_Plaintext(z_Plaintext),
    .Decryption_ready(Decryption_ready)
  );

  // Clock generation
  always #5 clk = ~clk;

  // Reset generation
  initial begin
    clk = 0;
    reset = 1;
    #10 reset = 0;
  end

  // Stimulus
  initial begin
    
    // plain text is P = ((X+1), (x+1)))
    x_C1  = 3'b111;
    y_C1 =  3'b000;
    z_C1 =  3'b110;
    x_C2 =  3'b100;
    y_C2 =  3'b101;
    z_C2 =  3'b110;


    #1000;
    // Add more test cases if needed

    $finish;
  end

endmodule
